library verilog;
use verilog.vl_types.all;
entity prod_tb is
end prod_tb;
