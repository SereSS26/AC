library verilog;
use verilog.vl_types.all;
entity patt_tb is
end patt_tb;
