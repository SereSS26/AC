library verilog;
use verilog.vl_types.all;
entity sm_unit_tb is
end sm_unit_tb;
