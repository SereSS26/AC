library verilog;
use verilog.vl_types.all;
entity mux_2s_tb is
    generic(
        W               : integer := 4
    );
end mux_2s_tb;
