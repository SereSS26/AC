library verilog;
use verilog.vl_types.all;
entity rot_r_tb is
end rot_r_tb;
