library verilog;
use verilog.vl_types.all;
entity div_by_6_tb is
end div_by_6_tb;
