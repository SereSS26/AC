library verilog;
use verilog.vl_types.all;
entity reg_parl_tb is
end reg_parl_tb;
