library verilog;
use verilog.vl_types.all;
entity minimization_tb is
end minimization_tb;
