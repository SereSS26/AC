library verilog;
use verilog.vl_types.all;
entity mul4_tb is
end mul4_tb;
