library verilog;
use verilog.vl_types.all;
entity comp_3b_tb is
end comp_3b_tb;
