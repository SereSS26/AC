library verilog;
use verilog.vl_types.all;
entity switch_tb is
end switch_tb;
