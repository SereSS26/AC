library verilog;
use verilog.vl_types.all;
entity tb_fsm_controller is
end tb_fsm_controller;
